module DCU();

endmodule